module mips(clk);
    input clk;
    reg[31:0] pc;
    wire[31:0] conba;
    
    
    
    
    
endmodule
